module reg_eg;
  reg y;
  wire a,b;
  initial begin
    y=a||b;
  end
endmodule
