module and_gate1(
    input a,
    input b,
    output y
    );
    assign y=a&b;
endmodule
