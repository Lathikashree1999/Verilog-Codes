module wire_eg;
  wire a,b,y;
  assign y = a&&b;
endmodule
